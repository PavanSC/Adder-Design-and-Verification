interface add_if(input bit clk);

parameter N=1;

logic  a;
 logic  b;
 logic c;
logic sum;
logic cout;
//logic rst;


endinterface



